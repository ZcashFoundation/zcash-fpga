module secp256k1_top (
  input                i_clk,
  input                i_rst,
  input                i_val,
  output logic         o_rdy,
  output logic         o_val
  
  
);

  
endmodule