module secp256k1_top ();
  
  
  // inversion
  
  // multiplication
  
  // addition
  
endmodule